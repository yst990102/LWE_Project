library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use work.configuration_set.all;

entity generate_dec is
    port (
        clk : in std_logic;

        q : in integer;
        s : in matrixS_1;
        RowU : in U_cell;
        RowV : in integer
        
        
    );
end generate_dec;

architecture Behavioral of generate_dec is

begin

end Behavioral;
